`include "digital_clock.v"

module tb();
    reg clk;
    reg rst;
    reg b;
    wire[3:0] hours_output;
    wire[6:0] minutes_output;
    wire[6:0] seconds_output;

    integer tb_iter;
    toplevel block(.clk(clk), .rst(rst), .b(b), .hours_output(hours_output), .minutes_output(minutes_output), .seconds_output(seconds_output));

    always
        #5 clk = ~clk;

    initial begin
        $dumpfile ("digital_clock.vcd");
        $dumpvars;

        clk = 0;
        rst = 0;
        block.hours_synth_0 = 0;
        block.hours_synth_1 = 0;
        block.hours_synth_2 = 0;
        block.hours_synth_3 = 0;
        block.minutes_synth_0 = 0;
        block.minutes_synth_1 = 0;
        block.minutes_synth_2 = 0;
        block.minutes_synth_3 = 0;
        block.minutes_synth_4 = 0;
        block.minutes_synth_5 = 0;
        block.minutes_synth_6 = 0;
        block.seconds_synth_0 = 0;
        block.seconds_synth_1 = 0;
        block.seconds_synth_2 = 0;
        block.seconds_synth_3 = 0;
        block.seconds_synth_4 = 0;
        block.seconds_synth_5 = 0;
        block.seconds_synth_6 = 0;
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        b = 1'd0;

        #10
        $finish;
    end
endmodule
